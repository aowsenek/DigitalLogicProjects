module Multiplexer(input [3:0]in0, input [3:0]in1, input [3:0]in2, input [3:0]in3, input [1:0] mode, output [3:0]o)
	assign o = in0;
endmodule