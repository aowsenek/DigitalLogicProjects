module Comparison(input [3:0]x, input [3:0]y, input [1:0] mode, output o);
	assign output = 1;
endmodule