module Arithmetic(input [7:0] i, input [1:0] mode, output [7:0] o);
	assign o = i;
endmodule