module Comparison(input [1:0] mode, input [3:0]x, input [3:0]y, output [3:0]o);
	assign o = x;
endmodule