module Project1_top(input [1:0]buttons, input [9:0]switches, output [9:0]LEDs, output [6:0]Hex1In, output [6:0]Hex2In);
//	SevenSegment Hex2(buttons, Hex1In[6:0]);
//	SevenSegment Hex1(switches[7:4], Hex2In[6:0]);
//	Logical test(switches[7:0], buttons, LEDs[7:0]);
endmodule 